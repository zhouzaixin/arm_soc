module cmsdk_top();



endmodule
